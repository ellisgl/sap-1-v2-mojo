`timescale 1ns / 1ps
module debounce(
    input      clk,
    input      in,
    output     out
);
	reg [19:0] ctr_d;
	reg [19:0] ctr_q;
	reg [1:0]  sync_d;
	reg [1:0]  sync_q;
 
	assign out = ctr_q == {20{1'b1}};
 
	always @(*)
	begin
		sync_d[0] = in;
		sync_d[1] = sync_q[0];
		ctr_d     = ctr_q + 1'b1;
 
		if (ctr_q == {20{1'b1}})
		begin
			ctr_d = ctr_q;
		end
 
		if (!sync_q[1])
		begin
			ctr_d = 20'd0;
		end
	end
 
	always @(posedge clk)
	begin
		ctr_q  <= ctr_d;
		sync_q <= sync_d;
	end
endmodule